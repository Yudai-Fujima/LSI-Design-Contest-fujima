library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity kernel_multiple is
  generic (
    CIN, COUT, HIN, WIN, K, S, P, HOUT, WOUT : integer;
    X_PLANE, Y_PLANE, DATA_WX, DATA_WW, ADDR_X_W, ADDR_W_W, ADDR_Y_W : integer
  );
  port (
    clk, rst, start : in std_logic;
    oc_sel : in integer;
    done : out std_logic;

    x_addr : out unsigned(ADDR_X_W-1 downto 0);
    x_dout : in  signed(DATA_WX-1 downto 0);

    w_raddr : out unsigned(ADDR_W_W-1 downto 0);
    w_dout  : in  signed(31 downto 0);

    y_raddr : out unsigned(ADDR_Y_W-1 downto 0);
    y_rdata : in  signed(31 downto 0);

    y_we    : out std_logic;
    y_waddr : out unsigned(ADDR_Y_W-1 downto 0);
    y_wdata : out signed(31 downto 0)
  );
end entity;

architecture rtl of kernel_multiple is

  component loop_counter
    generic (K, WIN, HIN, CIN : integer);
    port (
      clk, rst, step : in std_logic;
      kx, ky, ix, iy, ic : out integer;
      done : out std_logic
    );
  end component;

  component kernel_multiple_1
    generic (S, P, HOUT, WOUT, Y_PLANE, DATA_WIDTH : integer);
    port (
      iy, ix, ky, kx, ocv : in integer;
      x_in, w_in : in signed(DATA_WIDTH-1 downto 0);
      addr_y : out integer;
      prod_out : out signed(DATA_WIDTH-1 downto 0);
      valid : out std_logic
    );
  end component;

  component multiple
    generic (DATA_WIDTH : integer);
    port (
      x_in, w_in : in signed(DATA_WIDTH-1 downto 0);
      p_out : out signed(31 downto 0)
    );
  end component;

  component adder
    port (
      acc_in  : in signed(31 downto 0);
      prod_in : in signed(31 downto 0);
      sum_out : out signed(31 downto 0)
    );
  end component;

  type state_t is (
    IDLE,
    X_SETUP, X_WAIT, X_LATCH,
    W_SETUP, W_WAIT, W_LATCH,
    CALC_AND_READ_Y, WAIT_Y, ADD_WRITE,
    STEP_LOOP, POST_STEP,
    FINISH
  );
  signal st : state_t := IDLE;

  signal step_cnt  : std_logic := '0';
  signal loop_done : std_logic := '0';

  signal kx, ky, ix, iy, ic : integer := 0;

  signal x_reg, w_reg : signed(DATA_WX-1 downto 0) := (others=>'0');

  signal km1_addr_y     : integer := 0;
  signal km1_prod_dummy : signed(DATA_WX-1 downto 0) := (others=>'0');
  signal km1_valid      : std_logic := '0';

  signal mult_prod_32 : signed(31 downto 0) := (others=>'0');
  signal add_sum_32   : signed(31 downto 0) := (others=>'0');

  signal r_y_raddr_sig : unsigned(ADDR_Y_W-1 downto 0) := (others=>'0');
  signal cnt_rst       : std_logic;

  -- q(���b�`�������[�v�l)
  signal kx_q, ky_q, ix_q, iy_q, ic_q : integer := 0;

  -- ��prime����FOC���Ƃɍŏ���1�񂾂������Ȃ�
  signal priming : std_logic := '1';

  -- ��start�����オ�茟�o
  signal start_d    : std_logic := '0';
  signal start_rise : std_logic;
  -- �y�ǉ��z�o�C�g�I��p�̐M���i0�`3��ێ��j
  signal w_byte_sel : integer range 0 to 3 := 0;

begin

  -- loop_counter �� IDLE �̊Ԃ̓��Z�b�g
  --cnt_rst <= '1' when (rst = '1' or st = IDLE) else '0';
  cnt_rst <= '1' when (rst='1' or start_rise='1') else '0';

  u_counter : loop_counter
    generic map (K=>K, WIN=>WIN, HIN=>HIN, CIN=>CIN)
    port map (clk, cnt_rst, step_cnt, kx, ky, ix, iy, ic, loop_done);

  -- ��km1 �ɂ� q ������i���Ȃ��̍\���ێ��j
  u_km1 : kernel_multiple_1
    generic map (S=>S, P=>P, HOUT=>HOUT, WOUT=>WOUT, Y_PLANE=>Y_PLANE, DATA_WIDTH=>DATA_WX)
    port map (iy_q, ix_q, ky_q, kx_q, oc_sel, x_reg, w_reg, km1_addr_y, km1_prod_dummy, km1_valid);

  u_mult_32 : multiple
    generic map (DATA_WIDTH => DATA_WX)
    port map (x_reg, w_reg, mult_prod_32);

  u_adder_32 : adder
    port map (y_rdata, mult_prod_32, add_sum_32);

  y_raddr <= r_y_raddr_sig;
  y_wdata <= add_sum_32;

  -- ��start�����オ��
  start_rise <= start and (not start_d);

  process(clk, rst)
    variable widx : integer;
  begin
    if rst = '1' then
      st <= IDLE;

      step_cnt <= '0';
      done     <= '0';

      x_addr  <= (others=>'0');
      w_raddr <= (others=>'0');

      x_reg <= (others=>'0');
      w_reg <= (others=>'0');

      y_we    <= '0';
      y_waddr <= (others=>'0');

      r_y_raddr_sig <= (others=>'0');

      kx_q <= 0; ky_q <= 0; ix_q <= 0; iy_q <= 0; ic_q <= 0;

      priming <= '1';
      start_d <= '0';

    elsif rising_edge(clk) then
      -- -----------------------------------------
      -- start edge �̕ێ�
      -- -----------------------------------------
      start_d <= start;

      -- ���������́F
      -- start �������オ������u����OC�̍ŏ��͎̂Ă�v�ɖ߂�
      if start_rise = '1' then
        priming <= '1';
        -- q�������Ŋm���ɏ������i�ŏ��� addr �v�Z�����肳����j
        kx_q <= 0; ky_q <= 0; ix_q <= 0; iy_q <= 0; ic_q <= 0;
      end if;

      -- �f�t�H���g
      step_cnt <= '0';
      y_we     <= '0';
      done     <= '0';

      case st is
        when IDLE =>
          -- ��IDLE�ł� priming ��G��Ȃ��i�����d�v�j
          if start = '1' then
            st <= X_SETUP;
          end if;

        when X_SETUP =>
          x_addr <= to_unsigned(ic_q * X_PLANE + iy_q * WIN + ix_q, ADDR_X_W);
          st <= X_WAIT;

        when X_WAIT =>
          st <= X_LATCH;

        when X_LATCH =>
          x_reg <= x_dout;
          st <= W_SETUP;

        -- =========================================================
        -- �y�C���ӏ� 1�z �A�h���X�v�Z�ƃo�C�g�I���ʒu�̌���
        -- =========================================================
        when W_SETUP =>
          -- �{���̒ʂ��ԍ����v�Z
          widx := (ic_q * K + ky_q) * K + kx_q;
          
          -- RAM�A�h���X�� 1/4 (�����̊���Z�Ŏ����I�ɐ؂�̂�)
          w_raddr <= to_unsigned(widx / 4, ADDR_W_W);
          
          -- 32bit���̂ǂ̈ʒu�� (�]���ۑ�)
          w_byte_sel <= widx mod 4;
          
          st <= W_WAIT;

        when W_WAIT =>
          st <= W_LATCH;

        -- =========================================================
        -- �y�C���ӏ� 2�z �f�[�^�̐؂�o���E�����g���E2�{��(���V�t�g)
        -- =========================================================
        when W_LATCH =>
          -- w_dout(32bit)����8bit�؂�o�� -> DATA_WX(16bit��)�Ɋg�� -> 1�r�b�g���V�t�g(2�{)
          
          case w_byte_sel is
            when 0 => 
              -- Bits 7-0
              w_reg <= shift_left(resize(w_dout(7 downto 0), DATA_WX), 1);
            when 1 => 
              -- Bits 15-8
              w_reg <= shift_left(resize(w_dout(15 downto 8), DATA_WX), 1);
            when 2 => 
              -- Bits 23-16
              w_reg <= shift_left(resize(w_dout(23 downto 16), DATA_WX), 1);
            when 3 => 
              -- Bits 31-24
              w_reg <= shift_left(resize(w_dout(31 downto 24), DATA_WX), 1);
            when others =>
              w_reg <= (others => '0');
          end case;

          st <= CALC_AND_READ_Y;

        when CALC_AND_READ_Y =>
          if km1_valid = '1' and km1_addr_y >= 0 and km1_addr_y < (COUT * Y_PLANE) then
            r_y_raddr_sig <= to_unsigned(km1_addr_y, ADDR_Y_W);
            st <= WAIT_Y;
          else
            st <= STEP_LOOP;
          end if;

        when WAIT_Y =>
          st <= ADD_WRITE;

        when ADD_WRITE =>
          -- ��prime�FOC�ؑ֒���� "�ŏ���1��" �͏����Ȃ�
          if priming = '0' then
            y_we    <= '1';
            y_waddr <= r_y_raddr_sig;
          end if;

          -- ��������1��ڂ����������̂ŉ���
          priming <= '0';
          st <= STEP_LOOP;

        when STEP_LOOP =>
          step_cnt <= '1';
          st <= POST_STEP;

        when POST_STEP =>
          -- loop_counter �̍X�V�� q �ɔ��f
          kx_q <= kx; ky_q <= ky; ix_q <= ix; iy_q <= iy; ic_q <= ic;

          if loop_done = '1' then
            st <= FINISH;
          else
            st <= X_SETUP;
          end if;

        when FINISH =>
          done <= '1';
          if start = '0' then
            st <= IDLE;
          end if;

      end case;
    end if;
  end process;

end architecture;